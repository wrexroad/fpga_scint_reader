library verilog;
use verilog.vl_types.all;
entity NOT_1 is
    port(
        a               : in     vl_logic;
        not_a           : out    vl_logic
    );
end NOT_1;
